`resetall
`timescale 1ns / 1ps
// `default_nettype none


module ctrl_reg #(
  parameter        NUM_REGS    = 4,                              // liczba rejestrow
  parameter        REG_WIDTH   = 32,                             // szerokosc rejestrow (w bitach)
  parameter [31:0] IP_ADRESS   = {8'd192, 8'd168, 8'd1, 8'd128}, // adres IP komputera
  parameter [15:0] PORT_NUMBER = 16'd1234                        // numer portu
)(
  input  wire i_clk,
  input  wire i_rst,

  input  wire [7:0] i_rx_udp_payload_axis_tdata,
  input  wire       i_rx_udp_payload_axis_tvalid,
  input  wire       i_rx_udp_payload_axis_tlast,
  output wire       o_rx_udp_payload_axis_tready,

  output wire [7:0] o_tx_udp_payload_axis_tdata,
  output wire       o_tx_udp_payload_axis_tvalid,
  output wire       o_tx_udp_payload_axis_tlast,
  input  wire       i_tx_udp_payload_axis_tready,

  input  wire [15:0] i_port_nbr,
  input  wire [31:0] i_ip_adr,

  output wire [REG_WIDTH-1:0] o_reg_0,
  output wire [REG_WIDTH-1:0] o_reg_1,
  output wire [REG_WIDTH-1:0] o_reg_2,
  output wire [REG_WIDTH-1:0] o_reg_3
);


reg [REG_WIDTH-1:0] registers [0:NUM_REGS-1];

assign o_reg_0 = registers[0];
assign o_reg_1 = registers[1];
assign o_reg_2 = registers[2];
assign o_reg_3 = registers[3];

localparam [2:0] S_IDLE         = 3'd0;
localparam [2:0] S_WAIT_REG_NBR = 3'd1;
localparam [2:0] S_WAIT_CMD     = 3'd2;
localparam [2:0] S_WRITE_REG    = 3'd3;
localparam [2:0] S_READ_REG     = 3'd4;
localparam [2:0] S_ECHO         = 3'd5;

localparam [7:0] ASCII_NBR_BASE = 8'h30;
localparam [7:0] ASCII_W_UPPER  = 8'h57;
localparam [7:0] ASCII_W_LOWER  = 8'h77;
localparam [7:0] ASCII_R_UPPER  = 8'h52;
localparam [7:0] ASCII_R_LOWER  = 8'h72;
localparam [7:0] ASCII_COLON    = 8'h3A;

reg           [2:0] r_state, next_state;
reg           [2:0] r_reg_number, next_reg_number;
reg [REG_WIDTH-1:0] r_write_data, next_write_data;
reg           [4:0] r_write_byte_cnt, next_write_byte_cnt;
reg [REG_WIDTH-1:0] r_read_data, next_read_data;
reg           [2:0] r_read_byte_cnt, next_read_byte_cnt;
reg                 r_read_active, next_read_active;
reg                 r_rx_udp_payload_axis_tready;

reg           [7:0] r_tx_data;
reg                 r_tx_valid, next_tx_valid;
reg                 r_tx_last;
reg           [2:0] r_send_byte_cnt;

wire en;

integer i;
always @(posedge i_clk) begin
  if (i_rst) begin
    for (i = 0; i < NUM_REGS; i = i + 1) begin
      registers[i] <= 0;
    end
  end
end


assign en = (i_ip_adr==IP_ADRESS && i_port_nbr==PORT_NUMBER) ? 1'b1 : 1'b0;


always @(posedge i_clk)
begin: FSM_REGISTERS
  if (i_rst) begin
    r_state          <= S_IDLE;
    r_reg_number     <= 0;
    r_write_data     <= 0;
    r_write_byte_cnt <= 0;
    r_read_data      <= 0;
    r_read_byte_cnt  <= 0;
    r_read_active    <= 0;
  // end else begin
  end else if (en) begin
    r_state          <= next_state;
    r_reg_number     <= next_reg_number;
    r_write_data     <= next_write_data;
    r_write_byte_cnt <= next_write_byte_cnt;
    r_read_data      <= next_read_data;
    r_read_byte_cnt  <= next_read_byte_cnt;
    r_read_active    <= next_read_active;
  end
end // FSM_REGISTERS


always @(*)
begin: FSM_COMBINATIONAL
  next_state          = r_state;
  next_reg_number     = r_reg_number;
  next_write_data     = r_write_data;
  next_write_byte_cnt = r_write_byte_cnt;
  next_read_data      = r_read_data;
  next_read_byte_cnt  = r_read_byte_cnt;
  next_read_active    = r_read_active;
        next_tx_valid  = 0;

  case (r_state)
    S_IDLE: begin
      if (i_rx_udp_payload_axis_tvalid) begin
        if (i_rx_udp_payload_axis_tdata == ASCII_COLON) begin // czy odebrany znak to ':'?
          next_state          = S_WAIT_REG_NBR;
          next_write_byte_cnt = 0;
        end else begin // czy odebrany znak jest inny ni? ':'?
          next_state          = S_ECHO;
          next_tx_valid       = 1;
        end
      end
    end // S_IDLE

    S_WAIT_REG_NBR: begin
      if (i_rx_udp_payload_axis_tvalid) begin
        if (i_rx_udp_payload_axis_tdata >= ASCII_NBR_BASE &&
            i_rx_udp_payload_axis_tdata < (ASCII_NBR_BASE+NUM_REGS)) begin // czy numer rejestru jest w zakresie?
          next_state      = S_WAIT_CMD;
          next_reg_number = i_rx_udp_payload_axis_tdata - ASCII_NBR_BASE;
        end else begin // czy numer rejestru jest poza zakresem?
          next_state    = S_ECHO; // S_IDLE
          next_tx_valid = 1;
        end
      end
    end // S_WAIT_REG

    S_WAIT_CMD: begin
      if (i_rx_udp_payload_axis_tvalid) begin
        if (i_rx_udp_payload_axis_tdata == ASCII_W_UPPER ||
            i_rx_udp_payload_axis_tdata == ASCII_W_LOWER) begin // czy modyfiakcja zawartosci rejestru?
          next_state          = S_WRITE_REG;
          next_write_data     = 0;
          next_write_byte_cnt = 0;
        end else if (i_rx_udp_payload_axis_tdata == ASCII_R_UPPER ||
                     i_rx_udp_payload_axis_tdata == ASCII_R_LOWER) begin // czy odczyt z rejestru?
          next_state          = S_READ_REG;
          next_read_byte_cnt  = (REG_WIDTH/8)-1;
          next_read_data      = registers[r_reg_number];
          next_read_active    = 1;
        end else begin // czy komenda nieznana?
          next_state          = S_ECHO; // S_IDLE
          next_tx_valid       = 1;
        end
      end
    end // S_WAIT_CMD

    S_WRITE_REG: begin
      if (i_rx_udp_payload_axis_tvalid) begin
        next_write_data = (r_write_data << 8) | i_rx_udp_payload_axis_tdata;
        next_write_byte_cnt = r_write_byte_cnt + 1;
        if (r_write_byte_cnt < (REG_WIDTH/8) - 1) begin // czy jest w zakresie?
          if (i_rx_udp_payload_axis_tlast) begin // czy skonczyl odbierac?
            registers[r_reg_number] <= next_write_data;
            next_state              = S_IDLE;
          end
        end else begin // czy zapisano caly rejestr?
          next_state = S_IDLE;
          registers[r_reg_number] <= next_write_data;
        end
      end
    end // S_WRITE_REG

    S_READ_REG: begin
      if (r_read_active && i_tx_udp_payload_axis_tready) begin
        if (r_read_byte_cnt == 0) begin // czy wyslano cala zawartosc? 
          next_read_active   = 0;
          next_state         = S_IDLE;
        end else begin // czy kontynuowac wysylanie?
          next_read_byte_cnt = r_read_byte_cnt - 1;
        end
      end
    end // S_READ_REG

    S_ECHO: begin
      next_tx_valid   = 1;
      if (i_rx_udp_payload_axis_tvalid && i_rx_udp_payload_axis_tlast) begin
        next_state    = S_IDLE;
        next_tx_valid = 0;
      end
    end // S_ECHO
  endcase // state_reg
end // FSM_COMBINATIONAL


// wysylanie danych
always @(posedge i_clk) begin
  if (i_rst) begin
    r_tx_data       <= 0;
    r_tx_valid      <= 0;
    r_tx_last       <= 0;
    r_send_byte_cnt <= 0;

  // end else begin
  end else if (en) begin
    if (r_state == S_READ_REG && r_read_active) begin
      if (i_tx_udp_payload_axis_tready) begin
        case (r_read_byte_cnt) // wybierz odpowiedni bajt z rejestru do wyslania
          0: r_tx_data <= r_read_data[ 7: 0];
          1: r_tx_data <= r_read_data[15: 8];
          2: r_tx_data <= r_read_data[23:16];
          3: r_tx_data <= r_read_data[31:24];
          default: r_tx_data <= 0;
        endcase // r_read_byte_cnt
        r_tx_valid <= 1;
        if (r_read_byte_cnt == 0) begin
          r_tx_last <= 1;
        end
      end
    end else if (r_state == S_ECHO) begin
      if (i_rx_udp_payload_axis_tvalid) begin
        r_tx_data  <= i_rx_udp_payload_axis_tdata;
        r_tx_valid <= 1;
        r_tx_last  <= i_rx_udp_payload_axis_tlast;
      end
    end else begin
      r_tx_data  <= i_rx_udp_payload_axis_tdata;
      r_tx_valid <= next_tx_valid;
      r_tx_last  <= 0;
    end
  end
end


assign o_rx_udp_payload_axis_tready = (r_state == S_IDLE) || 
                                      (r_state == S_WAIT_REG_NBR) || 
                                      (r_state == S_WAIT_CMD) || 
                                      (r_state == S_WRITE_REG) || 
                                      (r_state == S_ECHO && i_tx_udp_payload_axis_tready);

assign o_tx_udp_payload_axis_tdata  = r_tx_data;
assign o_tx_udp_payload_axis_tvalid = r_tx_valid;
assign o_tx_udp_payload_axis_tlast  = r_tx_last;


endmodule // ctrl_reg